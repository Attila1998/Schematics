* C:\Users\pal.janos.attila\Desktop\Integ-4szog.sch

* Schematics Version 9.1 - Web Update 1
* Wed Oct 30 11:32:14 2019



** Analysis setup **
.tran 0ns 1s 0 0.1m
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Integ-4szog.net"
.INC "Integ-4szog.als"


.probe


.END
